module pc_register #(parameter width = 32)
(
    input clk,
    input load,
    input [width-1:0] in,
    output logic [width-1:0] out
);

logic [width-1:0] data;

/* Altera device registers are 0 at power on. Specify this
 * so that Modelsim works as expected.
 */
initial
begin
    data = 32'h00000060;
end

always_ff @(posedge clk)
begin
    if (load)
    begin
        data = in;
    end
	else /*DO NOTHING*/;
end

always_comb
begin
    out = data;
end

endmodule : pc_register
